interface intf();
  logic a,b,cin,sum,cout;
endinterface
