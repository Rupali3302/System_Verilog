interface intf();
  logic clock;
  logic reset;
  logic [4:0] in1;
  logic [4:0] in2; 
  logic [5:0] out; 
endinterface: intf
